module test();

wire a;
endmodule

