module test();


endmodule

