module test();

wire b,c;
endmodule

