module test();
//test20221215ㄝ, change2
wire b,c;
endmodule

