module test();

wire b;
endmodule

