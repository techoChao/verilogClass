module test();
//test20221215
wire b,c;
endmodule

